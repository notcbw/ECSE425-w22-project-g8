-- decode