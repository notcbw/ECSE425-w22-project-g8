-- memory