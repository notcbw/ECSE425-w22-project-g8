-- execute