-- put all components together