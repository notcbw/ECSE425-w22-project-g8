-- write back