-- fetch